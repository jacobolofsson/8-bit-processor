entity my_ram
end entity;