entity my_adress_register
end entity;