entity my_ALU
end entity;