entity my_control_unit
end entity;