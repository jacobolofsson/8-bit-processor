entity my_program_counter
end entity;