entity my_loop_counter
end entity;